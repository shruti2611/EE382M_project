interface mesi_output_interface();


endinterface : mesi_output_interface