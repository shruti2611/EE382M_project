interface mesi_input_interface(input clk, input rst);

endinterface : mesi_input_interface