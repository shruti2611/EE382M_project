class input_tx extends uvm_sequence_item;
	`uvm_object_utils(input_tx);

	//Specify inputs and constraints

	function new(string name);
		super.new(name);
	
	endfunction : newstring name

endclass : input_tx